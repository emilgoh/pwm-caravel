VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_pwm
  CLASS BLOCK ;
  FOREIGN user_proj_pwm ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2964.840 4.000 2965.440 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.880 4.000 366.480 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_in[14]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2764.920 4.000 2765.520 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2565.000 4.000 2565.600 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2365.080 4.000 2365.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2165.160 4.000 2165.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1965.240 4.000 1965.840 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1765.320 4.000 1765.920 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1565.400 4.000 1566.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1365.480 4.000 1366.080 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2831.560 4.000 2832.160 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END io_oeb[14]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2631.640 4.000 2632.240 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2431.720 4.000 2432.320 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2231.800 4.000 2232.400 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2031.880 4.000 2032.480 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1831.960 4.000 1832.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1632.040 4.000 1632.640 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1432.120 4.000 1432.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1232.200 4.000 1232.800 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1032.280 4.000 1032.880 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2898.200 4.000 2898.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_out[14]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2698.280 4.000 2698.880 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2498.360 4.000 2498.960 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2298.440 4.000 2299.040 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2098.520 4.000 2099.120 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1898.600 4.000 1899.200 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.680 4.000 1699.280 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 194.120 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 176.210 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 176.210 4.280 ;
      LAYER met3 ;
        RECT 3.990 2965.840 176.230 2986.725 ;
        RECT 4.400 2964.440 176.230 2965.840 ;
        RECT 3.990 2899.200 176.230 2964.440 ;
        RECT 4.400 2897.800 176.230 2899.200 ;
        RECT 3.990 2832.560 176.230 2897.800 ;
        RECT 4.400 2831.160 176.230 2832.560 ;
        RECT 3.990 2765.920 176.230 2831.160 ;
        RECT 4.400 2764.520 176.230 2765.920 ;
        RECT 3.990 2699.280 176.230 2764.520 ;
        RECT 4.400 2697.880 176.230 2699.280 ;
        RECT 3.990 2632.640 176.230 2697.880 ;
        RECT 4.400 2631.240 176.230 2632.640 ;
        RECT 3.990 2566.000 176.230 2631.240 ;
        RECT 4.400 2564.600 176.230 2566.000 ;
        RECT 3.990 2499.360 176.230 2564.600 ;
        RECT 4.400 2497.960 176.230 2499.360 ;
        RECT 3.990 2432.720 176.230 2497.960 ;
        RECT 4.400 2431.320 176.230 2432.720 ;
        RECT 3.990 2366.080 176.230 2431.320 ;
        RECT 4.400 2364.680 176.230 2366.080 ;
        RECT 3.990 2299.440 176.230 2364.680 ;
        RECT 4.400 2298.040 176.230 2299.440 ;
        RECT 3.990 2232.800 176.230 2298.040 ;
        RECT 4.400 2231.400 176.230 2232.800 ;
        RECT 3.990 2166.160 176.230 2231.400 ;
        RECT 4.400 2164.760 176.230 2166.160 ;
        RECT 3.990 2099.520 176.230 2164.760 ;
        RECT 4.400 2098.120 176.230 2099.520 ;
        RECT 3.990 2032.880 176.230 2098.120 ;
        RECT 4.400 2031.480 176.230 2032.880 ;
        RECT 3.990 1966.240 176.230 2031.480 ;
        RECT 4.400 1964.840 176.230 1966.240 ;
        RECT 3.990 1899.600 176.230 1964.840 ;
        RECT 4.400 1898.200 176.230 1899.600 ;
        RECT 3.990 1832.960 176.230 1898.200 ;
        RECT 4.400 1831.560 176.230 1832.960 ;
        RECT 3.990 1766.320 176.230 1831.560 ;
        RECT 4.400 1764.920 176.230 1766.320 ;
        RECT 3.990 1699.680 176.230 1764.920 ;
        RECT 4.400 1698.280 176.230 1699.680 ;
        RECT 3.990 1633.040 176.230 1698.280 ;
        RECT 4.400 1631.640 176.230 1633.040 ;
        RECT 3.990 1566.400 176.230 1631.640 ;
        RECT 4.400 1565.000 176.230 1566.400 ;
        RECT 3.990 1499.760 176.230 1565.000 ;
        RECT 4.400 1498.360 176.230 1499.760 ;
        RECT 3.990 1433.120 176.230 1498.360 ;
        RECT 4.400 1431.720 176.230 1433.120 ;
        RECT 3.990 1366.480 176.230 1431.720 ;
        RECT 4.400 1365.080 176.230 1366.480 ;
        RECT 3.990 1299.840 176.230 1365.080 ;
        RECT 4.400 1298.440 176.230 1299.840 ;
        RECT 3.990 1233.200 176.230 1298.440 ;
        RECT 4.400 1231.800 176.230 1233.200 ;
        RECT 3.990 1166.560 176.230 1231.800 ;
        RECT 4.400 1165.160 176.230 1166.560 ;
        RECT 3.990 1099.920 176.230 1165.160 ;
        RECT 4.400 1098.520 176.230 1099.920 ;
        RECT 3.990 1033.280 176.230 1098.520 ;
        RECT 4.400 1031.880 176.230 1033.280 ;
        RECT 3.990 966.640 176.230 1031.880 ;
        RECT 4.400 965.240 176.230 966.640 ;
        RECT 3.990 900.000 176.230 965.240 ;
        RECT 4.400 898.600 176.230 900.000 ;
        RECT 3.990 833.360 176.230 898.600 ;
        RECT 4.400 831.960 176.230 833.360 ;
        RECT 3.990 766.720 176.230 831.960 ;
        RECT 4.400 765.320 176.230 766.720 ;
        RECT 3.990 700.080 176.230 765.320 ;
        RECT 4.400 698.680 176.230 700.080 ;
        RECT 3.990 633.440 176.230 698.680 ;
        RECT 4.400 632.040 176.230 633.440 ;
        RECT 3.990 566.800 176.230 632.040 ;
        RECT 4.400 565.400 176.230 566.800 ;
        RECT 3.990 500.160 176.230 565.400 ;
        RECT 4.400 498.760 176.230 500.160 ;
        RECT 3.990 433.520 176.230 498.760 ;
        RECT 4.400 432.120 176.230 433.520 ;
        RECT 3.990 366.880 176.230 432.120 ;
        RECT 4.400 365.480 176.230 366.880 ;
        RECT 3.990 300.240 176.230 365.480 ;
        RECT 4.400 298.840 176.230 300.240 ;
        RECT 3.990 233.600 176.230 298.840 ;
        RECT 4.400 232.200 176.230 233.600 ;
        RECT 3.990 166.960 176.230 232.200 ;
        RECT 4.400 165.560 176.230 166.960 ;
        RECT 3.990 100.320 176.230 165.560 ;
        RECT 4.400 98.920 176.230 100.320 ;
        RECT 3.990 33.680 176.230 98.920 ;
        RECT 4.400 32.280 176.230 33.680 ;
        RECT 3.990 10.715 176.230 32.280 ;
      LAYER met4 ;
        RECT 9.495 1564.855 19.025 2767.425 ;
  END
END user_proj_pwm
END LIBRARY

